module Clocked_
